module labka12(x, out);
input [3:0] x;
output out;



/*my_mux multiplexer(.data15(0), .data14(1), .data13(0), .data12(0),
					.data11(1), .data10(1),	.data9(0), .data8(0),
					.data7(0), .data6(0), .data5(1), .data4(0),
					.data3(1), .data2(1), .data1(1), .data0(0),
					.sel(x), .result(out));	*/
endmodule