library verilog;
use verilog.vl_types.all;
entity labka12 is
    port(
        x               : in     vl_logic_vector(3 downto 0);
        \out\           : out    vl_logic
    );
end labka12;
